`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:49:21 03/21/2024 
// Design Name: 
// Module Name:    prygen 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module prygen(X, Y, Z, Result);
    input X;
    input Y;
    input Z;
    output Result;
	 assign Result=X^Y^Z;
	 
endmodule
